--
--
--
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PI_controle is
    port();
end entity;

architecture main of PI_contorle is
begin
end architecture;