--
--
-- Author: Erick S. Dias
-- Last update: 26/03/25 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;